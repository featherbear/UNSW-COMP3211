-- Test communication between two ASIPs

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity test_network is
--  Port ( );
end test_network;

architecture Behavioural of test_network is

begin


end Behavioural;
